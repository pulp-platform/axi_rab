`include "BramPort.sv"

module axi4_bram_logger

  // Parameters {{{
  #(
    parameter AXI_ADDR_WIDTH  = 32,
    parameter AXI_ID_WIDTH    = 8,
    parameter AXI_LEN_WIDTH   = 8,
    parameter TIMESTAMP_WIDTH = 32,
    parameter BRAM_DATA_WIDTH = 32,
    parameter BRAM_ADDR_WIDTH = 18,
    parameter NUM_BRAMS       = 32
  )
  // }}}

  // Ports {{{
  (
    input  logic                                  Clk_CI,
    input  logic                                  Rst_RBI,

    // AXI Input
    input  logic                                  AxiValid_SI,
    input  logic  [AXI_ID_WIDTH-1:0]              AxiId_DI,
    input  logic  [AXI_ADDR_WIDTH-1:0]            AxiAddr_DI,
    input  logic  [AXI_LEN_WIDTH-1:0]             AxiLen_DI,

    // Control Input
    input  logic                                  Clear_SI,

    // Status Output
    output logic                                  Full_SO,

    // Interface to Internal BRAM
    // TODO: instantiate this interface with BRAM_ADDR_WIDTH and BRAM_DATA_WIDTH
    //BramPort #(
    //  .DATA_WIDTH(BRAM_ADDR_WIDTH),
    //  .ADDR_WIDTH(BRAM_ADDR_WIDTH))               Bram
    BramPort.Slave                                  Bram_PS
    // TODO, deprecated if the above works:
    //input  logic                                  BramClk_CI,
    //input  logic                                  BramRst_RI,
    //input  logic                                  BramEn_SI,
    //input  logic  [BRAM_ADDR_WIDTH-1:0]           BramAddr_SI,
    //output logic  [BRAM_DATA_WIDTH-1:0]           BramRd_DO,
    //input  logic  [BRAM_DATA_WIDTH-1:0]           BramWr_DI,
    //input  logic  [`log2(BRAM_DATA_WIDTH/4)-1:0]  BramWrEn_SI
  );
  // }}}

  // Signal Declarations {{{
  logic                                           Rst_R;

  logic                   [BRAM_DATA_WIDTH-1:0]   BramAWr_D;
  logic                   [16-1:0]                BramAAddr_S;
  logic [NUM_BRAMS-1:0]                           BramAWrEn_S;
  logic [NUM_BRAMS-1:0]   [BRAM_DATA_WIDTH-1:0]   BramBRd_D;
  logic [NUM_BRAMS-1:0]                           BramBWrEn_S;

  logic                                           BramAWr_S;
  // }}}

  // Register Declarations {{{
  reg [AXI_ADDR_WIDTH-1:0]        AxiAddr_DP,       AxiAddr_DN;
  reg [AXI_ID_WIDTH-1:0]          AxiId_DP,         AxiId_DN;
  reg [AXI_LEN_WIDTH-1:0]         AxiLen_DP,        AxiLen_DN;
  reg                             Full_SP,          Full_SN;
  reg [TIMESTAMP_WIDTH-1:0]       Timestamp_SP,     Timestamp_SN;
  reg [15:0]                      WrAddrCnt_SP,     WrAddrCnt_SN;

  enum {IDLE, WRITE_ADDR, WRITE_META}
                                  State_SP,         State_SN;
  // }}}

  assign Rst_R = ~Rst_RBI; // TODO: is the polarity of this reset suitable for the BRAM?

  // BRAM Instantiation and Port Assignment {{{
  genvar i;
  for (i = 0; i < NUM_BRAMS; i++) begin

    // RAMB36E1 {{{
    // RAMB36E1: 36K-bit Configurable Synchronous Block RAM
    //           Virtex-7
    // Xilinx HDL Language Template, version 2015.1
    RAMB36E1 #(
      // Address Collision Mode: "PERFORMANCE" or "DELAYED_WRITE"
      .RDADDR_COLLISION_HWCONFIG("DELAYED_WRITE"),
      // Collision check: Values ("ALL", "WARNING_ONLY", "GENERATE_X_ONLY" or "NONE")
      .SIM_COLLISION_CHECK("ALL"),
      // DOA_REG, DOB_REG: Optional output register (0 or 1)
      .DOA_REG(0),
      .DOB_REG(0),
      .EN_ECC_READ("FALSE"),                                                            // Enable ECC decoder,
                                                                                        // FALSE, TRUE
      .EN_ECC_WRITE("FALSE"),                                                           // Enable ECC encoder,
                                                                                        // FALSE, TRUE
      // INITP_00 to INITP_0F: Initial contents of the parity memory array
      .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
      // INIT_00 to INIT_7F: Initial contents of the data memory array
      .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_40(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_41(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_42(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_43(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_44(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_45(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_46(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_47(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_48(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_49(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_4A(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_4B(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_4C(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_4D(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_4E(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_4F(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_50(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_51(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_52(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_53(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_54(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_55(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_56(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_57(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_58(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_59(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_5A(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_5B(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_5C(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_5D(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_5E(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_5F(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_60(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_61(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_62(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_63(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_64(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_65(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_66(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_67(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_68(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_69(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_6A(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_6B(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_6C(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_6D(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_6E(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_6F(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_70(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_71(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_72(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_73(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_74(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_75(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_76(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_77(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_78(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_79(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_7A(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_7B(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_7C(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_7D(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_7E(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_7F(256'h0000000000000000000000000000000000000000000000000000000000000000),
      // INIT_A, INIT_B: Initial values on output ports
      .INIT_A(36'h000000000),
      .INIT_B(36'h000000000),
      // Initialization File: RAM initialization file
      .INIT_FILE("NONE"),
      // RAM Mode: "SDP" or "TDP"
      .RAM_MODE("TDP"),
      // RAM_EXTENSION_A, RAM_EXTENSION_B: Selects cascade mode ("UPPER", "LOWER", or "NONE")
      .RAM_EXTENSION_A("NONE"),
      .RAM_EXTENSION_B("NONE"),
      // READ_WIDTH_A/B, WRITE_WIDTH_A/B: Read/write width per port
      .READ_WIDTH_A(32),                                                                 // 0-72
      .READ_WIDTH_B(32),                                                                 // 0-36
      .WRITE_WIDTH_A(32),                                                                // 0-36
      .WRITE_WIDTH_B(32),                                                                // 0-72
      // RSTREG_PRIORITY_A, RSTREG_PRIORITY_B: Reset or enable priority ("RSTREG" or "REGCE")
      .RSTREG_PRIORITY_A("RSTREG"),
      .RSTREG_PRIORITY_B("RSTREG"),
      // SRVAL_A, SRVAL_B: Set/reset value for output
      .SRVAL_A(36'h000000000),
      .SRVAL_B(36'h000000000),
      // Simulation Device: Must be set to "7SERIES" for simulation behavior
      .SIM_DEVICE("7SERIES"),
      // WriteMode: Value on output upon a write ("WRITE_FIRST", "READ_FIRST", or "NO_CHANGE")
      .WRITE_MODE_A("WRITE_FIRST"),
      .WRITE_MODE_B("WRITE_FIRST")
    )
    // }}}

    // RAMB36E1_inst {{{
    RAMB36E1_inst (
      // Cascade Signals: 1-bit (each) output: BRAM cascade ports (to create 64kx1)
      .CASCADEOUTA(),     // 1-bit output: A port cascade
      .CASCADEOUTB(),     // 1-bit output: B port cascade
      // ECC Signals: 1-bit (each) output: Error Correction Circuitry ports
      .DBITERR(),             // 1-bit output: Double bit error status
      .ECCPARITY(),         // 8-bit output: Generated error correction parity
      .RDADDRECC(),         // 9-bit output: ECC read address
      .SBITERR(),             // 1-bit output: Single bit error status
      // Port A Data: 32-bit (each) output: Port A data
      .DOADO(),                 // 32-bit output: A port data/LSB data
      .DOPADOP(),             // 4-bit output: A port parity/LSB parity
      // Port B Data: 32-bit (each) output: Port B data
      .DOBDO(BramBRd_D[i]),                 // 32-bit output: B port data/MSB data
      .DOPBDOP(),             // 4-bit output: B port parity/MSB parity
      // Cascade Signals: 1-bit (each) input: BRAM cascade ports (to create 64kx1)
      .CASCADEINA(1'b0),       // 1-bit input: A port cascade
      .CASCADEINB(1'b0),       // 1-bit input: B port cascade
      // ECC Signals: 1-bit (each) input: Error Correction Circuitry ports
      .INJECTDBITERR(1'b0), // 1-bit input: Inject a double bit error
      .INJECTSBITERR(1'b0), // 1-bit input: Inject a single bit error
      // Port A Address/Control Signals: 16-bit (each) input: Port A address and control signals (read port
      // when RAM_MODE="SDP")
      .ADDRARDADDR(BramAAddr_S),     // 16-bit input: A port address/Read address
      .CLKARDCLK(Clk_CI),         // 1-bit input: A port clock/Read clock
      .ENARDEN(1'b1),             // 1-bit input: A port enable/Read enable
      .REGCEAREGCE(1'b1),     // 1-bit input: A port register enable/Register enable
      .RSTRAMARSTRAM(Rst_R), // 1-bit input: A port set/reset
      .RSTREGARSTREG(Rst_R), // 1-bit input: A port register set/reset
      .WEA(BramAWrEn_S[i]),                     // 4-bit input: A port write enable
      // Port A Data: 32-bit (each) input: Port A data
      .DIADI(BramAWr_D),                 // 32-bit input: A port data/LSB data
      .DIPADIP(4'b0000),             // 4-bit input: A port parity/LSB parity
      // Port B Address/Control Signals: 16-bit (each) input: Port B address and control signals (write port
      // when RAM_MODE="SDP")
      .ADDRBWRADDR(Bram_PS.Addr_S[12:0]),     // 16-bit input: B port address/Write address
      .CLKBWRCLK(Bram_PS.Clk_C),         // 1-bit input: B port clock/Write clock
      .ENBWREN(Bram_PS.En_S),             // 1-bit input: B port enable/Write enable
      .REGCEB(1'b1),               // 1-bit input: B port register enable
      .RSTRAMB(Bram_PS.Rst_R),             // 1-bit input: B port set/reset
      .RSTREGB(Bram_PS.Rst_R),             // 1-bit input: B port register set/reset
      .WEBWE(BramBWrEn_S[i]),                 // 8-bit input: B port write enable/Write enable
      // Port B Data: 32-bit (each) input: Port B data
      .DIBDI(Bram_PS.Wr_D),                 // 32-bit input: B port data/MSB data
      .DIPBDIP(4'b0000)              // 4-bit input: B port parity/MSB parity
    );
    // }}}

    // Port A Address-Dependent Write Enable {{{
    always_comb begin
      BramAWrEn_S[i] = '{default: '0};
      if (WrAddrCnt_SP[15:11] == i && BramAWr_S) begin
        BramAWrEn_S[i] = '{default: '1};
      end
    end
    // }}}

    // Port B Address-Dependent Write Enable {{{
    always_comb begin
      BramBWrEn_S[i] = '{default: '0};
      if (Bram_PS.Addr_S[17:13] == i) begin
        BramBWrEn_S[i] = Bram_PS.WrEn_S;
      end
    end
    // }}}

  end
  // }}}

  // Control FSM {{{
  always_comb
  begin
    // Default Assignments
    AxiAddr_DN  = AxiAddr_DP;
    AxiId_DN    = AxiId_DP;
    AxiLen_DN   = AxiLen_DP;
    BramAWr_D   = 0;
    BramAWr_S   = 0;
    State_SN    = State_SP;

    // Log AXI transfers if BRAM is not full.
    if (~Full_SP) begin
      case (State_SP)
        IDLE: begin
          if (AxiValid_SI) begin
            // Write timestamp to BRAM.
            BramAWr_D   = Timestamp_SP;
            BramAWr_S   = 1;

            // Latch AXI data.
            AxiAddr_DN  = AxiAddr_DI;
            AxiId_DN    = AxiId_DI;
            AxiLen_DN   = AxiLen_DI;

            State_SN    = WRITE_ADDR;
          end
        end
        WRITE_ADDR: begin
          // Write AXI address to BRAM.
          BramAWr_D = AxiAddr_DP;
          BramAWr_S = 1;

          State_SN  = WRITE_META;
        end
        WRITE_META: begin
          // Write AXI metadata to BRAM.
          BramAWr_D = {AxiId_DP, AxiLen_DP};
          BramAWr_S = 1;

          State_SN  = IDLE;
        end
      endcase
    end
  end
  // }}}

  // BRAM Write Address Generation {{{
  assign BramAAddr_S = WrAddrCnt_SP[10:0] << 2;
  always_comb
  begin
    WrAddrCnt_SN  = WrAddrCnt_SP;
    if (BramAWr_S) begin
      WrAddrCnt_SN = WrAddrCnt_SP + 1;
      if (WrAddrCnt_SP == $high(WrAddrCnt_SP)) begin
        WrAddrCnt_SN  = 0;
      end
    end
  end
  // }}}

  // BRAM Full Handler {{{
  always_comb
  begin
    Full_SN = Full_SP;
    if (WrAddrCnt_SP == $high(WrAddrCnt_SP)) begin
      Full_SN = 1;
    end
    // TODO: clearing
  end
  // }}}

  // Timestamp Counter {{{
  always_comb
  begin
    Timestamp_SN = Timestamp_SP + 1;
    if (Timestamp_SP == $high(Timestamp_SP)) begin
      Timestamp_SN = 0;
    end
  end
  // }}}

  // Flip-Flops {{{
  always_ff @ (posedge Clk_CI)
  begin
    if (~Rst_RBI) begin
      AxiAddr_DP    <= 0;
      AxiId_DP      <= 0;
      AxiLen_DP     <= 0;
      Full_SP       <= 0;
      Timestamp_SP  <= 0;
      WrAddrCnt_SP  <= 0;
    end else begin
      AxiAddr_DP    <= AxiAddr_DN;
      AxiId_DP      <= AxiId_DN;
      AxiLen_DP     <= AxiLen_DN;
      Full_SP       <= Full_SN;
      Timestamp_SP  <= Timestamp_SN;
      WrAddrCnt_SP  <= WrAddrCnt_SN;
    end
  end
  // }}}

  // BRAM Output Port Multiplexer
  assign Bram_PS.Rd_D = BramBRd_D[Bram_PS.Addr_S[17:13]];

  assign Full_SO = Full_SP;

endmodule

// vim: ts=2 sw=2 sts=2 et nosmartindent autoindent foldmethod=marker
