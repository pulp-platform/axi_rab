/* Copyright (C) 2017 ETH Zurich, University of Bologna
 * All rights reserved.
 *
 * This code is under development and not yet released to the public.
 * Until it is released, the code is under the copyright of ETH Zurich and
 * the University of Bologna, and may contain confidential and/or unpublished
 * work. Any reuse/redistribution is strictly forbidden without written
 * permission from ETH Zurich.
 *
 * Bug fixes and contributions will eventually be released under the
 * SolderPad open hardware license in the context of the PULP platform
 * (http://www.pulp-platform.org), under the copyright of ETH Zurich and the
 * University of Bologna.
 */

`include "ulpsoc_defines.sv"

//`define TLB_MULTIHIT

import CfMath::log2;

time clk_period = 10ns;    // clock generated by ARM

task tb_wait(input int cycles);
   #(clk_period*cycles);
endtask // tb_wait

module rab_tb
 #(
   parameter C_AXI_DATA_WIDTH    = 64,
   parameter C_AXICFG_DATA_WIDTH = 32,
   parameter C_AXI_ID_WIDTH      = 8,
   parameter C_AXI_USER_WIDTH    = 6,
   parameter BUFFER_SIZE = 8,
   parameter SRC_ID = 8,
   parameter TEST_NAME = "reg_rd_wr"
  )
;

   timeunit      1ps;
   timeprecision 1ps;

   localparam BUFFER_ADDR_BITS = log2(BUFFER_SIZE-1);
   localparam AXI_EXT_ADDR_WIDTH = 32;
   localparam MEM_ADDR_WIDTH     = AXI_EXT_ADDR_WIDTH-log2(C_AXI_DATA_WIDTH/8);

   logic   clk_i;         // input
   logic   rst_ni;      // input

   ///////////////////////////
   //
   // DUT - axi_rab_wrap
   //
   ///////////////////////////

   AXI_BUS #(
             .AXI_ADDR_WIDTH    ( 32                 ),
             .AXI_DATA_WIDTH    ( C_AXI_DATA_WIDTH   ),
             .AXI_ID_WIDTH      ( C_AXI_ID_WIDTH     ),
             .AXI_USER_WIDTH    ( C_AXI_USER_WIDTH   )
             ) tgen2rab();

   AXI_BUS #(
             .AXI_ADDR_WIDTH    ( AXI_EXT_ADDR_WIDTH ),
             .AXI_DATA_WIDTH    ( C_AXI_DATA_WIDTH   ),
             .AXI_ID_WIDTH      ( C_AXI_ID_WIDTH     ),
             .AXI_USER_WIDTH    ( C_AXI_USER_WIDTH   )
             ) rab2mem();

    AXI_BUS #(
             .AXI_ADDR_WIDTH    ( AXI_EXT_ADDR_WIDTH ),
             .AXI_DATA_WIDTH    ( C_AXI_DATA_WIDTH   ),
             .AXI_ID_WIDTH      ( C_AXI_ID_WIDTH     ),
             .AXI_USER_WIDTH    ( C_AXI_USER_WIDTH   )
             ) acp2mem();

    AXI_BUS #(
             .AXI_ADDR_WIDTH    ( 32                  ),
             .AXI_DATA_WIDTH    ( C_AXI_DATA_WIDTH    ),
             .AXI_ID_WIDTH      ( C_AXI_ID_WIDTH      ),
             .AXI_USER_WIDTH    ( C_AXI_USER_WIDTH    )
             ) rab_to_socbus_dummy();

    AXI_BUS #(
             .AXI_ADDR_WIDTH    ( 32                  ),
             .AXI_DATA_WIDTH    ( C_AXI_DATA_WIDTH    ),
             .AXI_ID_WIDTH      ( C_AXI_ID_WIDTH      ),
             .AXI_USER_WIDTH    ( C_AXI_USER_WIDTH    )
             ) rab_slave_dummy();


   logic          tgen2rab_eoc;
   logic          tgen2rab_fetch_en;
   logic [31:0]   tgen2rab_PASS;
   logic [31:0]   tgen2rab_FAIL;


   AXI_LITE #(
    .AXI_ADDR_WIDTH ( 32 ),
    .AXI_DATA_WIDTH ( C_AXICFG_DATA_WIDTH )
    ) rab_lite();

   logic        intr_mhf_full_o;
   logic        intr_miss_o;
   logic        intr_multi_o;
   logic        intr_prot_o;

   UNICAD_MEM_BUS_64 mem_if();
   UNICAD_MEM_BUS_64 mem_if_acp();


   axi_rab_wrap
   #(
      .N_SLICES               ( 32                 ),
      .AXI_EXT_ADDR_WIDTH     ( AXI_EXT_ADDR_WIDTH ),
      .AXI_ADDR_WIDTH         ( 32                 ),
      .AXI_DATA_WIDTH         ( C_AXI_DATA_WIDTH   ),
      .AXI_USER_WIDTH         ( C_AXI_USER_WIDTH   ),
      .AXI_LITE_ADDR_WIDTH    ( 32                 ),
      .AXI_LITE_DATA_WIDTH    ( 32                 ),
      .AXI_ID_EXT_S_WIDTH     ( C_AXI_ID_WIDTH     ),
      .AXI_ID_EXT_S_ACP_WIDTH ( C_AXI_ID_WIDTH     ),
      .AXI_ID_EXT_M_WIDTH     ( C_AXI_ID_WIDTH     ),
      .AXI_ID_SOC_S_WIDTH     ( C_AXI_ID_WIDTH     ),
      .AXI_ID_SOC_M_WIDTH     ( C_AXI_ID_WIDTH     ),
      .N_PORTS                ( 1                  )
     )
   DUT
     (
      .clk_i           ( clk_i               ),
      .rst_ni          ( rst_ni              ),

      .rab_to_socbus   ( rab_to_socbus_dummy ),
      .socbus_to_rab   ( tgen2rab            ),

      .rab_master      ( rab2mem             ),
      .rab_acp         ( acp2mem             ),
      .rab_slave       ( rab_slave_dummy     ),

      .rab_lite        ( rab_lite            ),

      .intr_miss_o     ( intr_miss_o         ),
      .intr_multi_o    ( intr_multi_o        ),
      .intr_prot_o     ( intr_prot_o         ),
      .intr_mhf_full_o ( intr_mhf_full_o     )
    );

   ///////////////////////////
   //
   // axi4lite verification ip
   //
   ///////////////////////////
   axi4lite_m_if axi4lite_m_if_0(clk_i);

   // Master write address channel
   assign rab_lite.aw_addr   = axi4lite_m_if_0.awaddr ;
   assign rab_lite.aw_valid  = axi4lite_m_if_0.awvalid;
   assign axi4lite_m_if_0.awready = rab_lite.aw_ready ;
   // Master write data channel
   assign rab_lite.w_data    = axi4lite_m_if_0.wdata  ;
   assign rab_lite.w_strb    = axi4lite_m_if_0.wstrb  ;
   assign rab_lite.w_valid   = axi4lite_m_if_0.wvalid ;
   assign axi4lite_m_if_0.wready  = rab_lite.w_ready  ;
   // Master write response channel
   assign axi4lite_m_if_0.bresp   = rab_lite.b_resp   ;
   assign axi4lite_m_if_0.bvalid  = rab_lite.b_valid  ;
   assign rab_lite.b_ready   = axi4lite_m_if_0.bready ;
   // Master read address channel
   assign rab_lite.ar_addr   = axi4lite_m_if_0.araddr ;
   assign rab_lite.ar_valid  = axi4lite_m_if_0.arvalid;
   assign axi4lite_m_if_0.arready = rab_lite.ar_ready ;
   // Master read data channel
   assign axi4lite_m_if_0.rdata   = rab_lite.r_data   ;
   assign axi4lite_m_if_0.rresp   = rab_lite.r_resp   ;
   assign axi4lite_m_if_0.rvalid  = rab_lite.r_valid  ;
   assign rab_lite.r_ready   = axi4lite_m_if_0.rready ;


  ///////////////////////////
  //
  // AXI TGEN Interface
  //
  ///////////////////////////
  TGEN_wrap
  #(
    .AXI4_ADDRESS_WIDTH ( 32               ),
    .AXI4_RDATA_WIDTH   ( C_AXI_DATA_WIDTH ),
    .AXI4_WDATA_WIDTH   ( C_AXI_DATA_WIDTH ),
    .AXI4_ID_WIDTH      ( C_AXI_ID_WIDTH   ),
    .AXI4_USER_WIDTH    ( C_AXI_USER_WIDTH ),
    .SRC_ID             ( SRC_ID           )
  )
  axi_m_if_0(
    .clk             ( clk_i             ),
    .rst_n           ( rst_ni            ),
    .axi_port_master ( tgen2rab          ),
    .eoc_o           ( tgen2rab_eoc      ),
    .fetch_en_i      ( tgen2rab_fetch_en ),
    .PASS_o          ( tgen2rab_PASS     ),
    .FAIL_o          ( tgen2rab_FAIL     )
  );

  ///////////////////////////
  //
  // Memory Interface
  //
  ///////////////////////////
  axi_mem_if_wrap
  #(
   .AXI_ADDRESS_WIDTH ( AXI_EXT_ADDR_WIDTH ),
   .AXI_DATA_WIDTH    ( C_AXI_DATA_WIDTH   ),
   .AXI_ID_WIDTH      ( C_AXI_ID_WIDTH     ),
   .AXI_USER_WIDTH    ( C_AXI_USER_WIDTH   )
  )
  axi_mem_if_0
  (
    .clk_i      ( clk_i   ),
    .rst_ni     ( rst_ni  ),
    .test_en_i  ( 1'b0    ),
    .axi_slave  ( rab2mem ),
    .mem_master ( mem_if  )
  );

  axi_mem_if_wrap
  #(
    .AXI_ADDRESS_WIDTH ( AXI_EXT_ADDR_WIDTH ),
    .AXI_DATA_WIDTH    ( C_AXI_DATA_WIDTH   ),
    .AXI_ID_WIDTH      ( C_AXI_ID_WIDTH     ),
    .AXI_USER_WIDTH    ( C_AXI_USER_WIDTH   )
  )
  axi_mem_if_acp
  (
    .clk_i      ( clk_i      ),
    .rst_ni     ( rst_ni     ),
    .test_en_i  ( 1'b0       ),
    .axi_slave  ( acp2mem    ),
    .mem_master ( mem_if_acp )
  );

  l2_ram
  #(
    .MEM_ADDR_WIDTH ( MEM_ADDR_WIDTH )
   )
  ram_0
  (
    .clk_i     ( clk_i  ),
    .rst_ni    ( rst_ni ),
    .mem_slave ( mem_if ),
    .test_en_i ( 1'b0   )
  );

  l2_ram
  #(
    .MEM_ADDR_WIDTH ( MEM_ADDR_WIDTH )
  )
  ram_0_acp
  (
    .clk_i     ( clk_i      ),
    .rst_ni    ( rst_ni     ),
    .mem_slave ( mem_if_acp ),
    .test_en_i ( 1'b0       )
  );

   ///////////////////////////
   //
   // Clock and Reset
   //
   ///////////////////////////
   initial
     begin
        rst_ni = 1'b1;
        tb_wait(1);
        rst_ni = 1'b0;
        tb_wait(10);
        rst_ni = 1'b1; // release reset
        tb_wait(10);
     end
   initial
     begin : clk_gen
        clk_i = 1'b1;
        #(clk_period/2-1);
        forever #(clk_period/2) clk_i = ~clk_i;
     end


  ///////////////////////////
  //
  //// Test
  //
  ///////////////////////////
  test
  #(
   .TEST_NAME ( TEST_NAME )
  )
  u_test();



   ///////////////////////////
   //
   ////  Monitors / Checkers
   //
   ///////////////////////////

   ////////////////////////////////////////////////////////////////////////////////////////
   /////////////////////////// Check axi_lite transactions ////////////////////////////////
   ////////////////////////////////////////////////////////////////////////////////////////
   bit [31:0] regblock[383:0], va_block[1023:0], pa_block[1023:0];
   int       unsigned regblock_w_addr,regblock_r_addr, ram_addr;
   int       unsigned error_num,error_miss=0,error_axi = 0, error_buf=0;

   //////// RAB Registers

   // Write data into reg model
   always_comb begin
      if (rab_lite.aw_valid == 1 && rab_lite.aw_addr < 32'h4000) begin
         regblock_w_addr = rab_lite.aw_addr;
      end

      if (rab_lite.w_valid == 1 && rab_lite.aw_addr < 32'h4000) begin
         regblock[regblock_w_addr/4] =  rab_lite.w_data;
         $display("Register Write detected at monitor. Address = %h",regblock_w_addr);
      end
   end // always_comb begin

   // Check if read data is correct in reg model
   always_comb begin
      if (rab_lite.ar_valid == 1 && rab_lite.ar_addr < 32'h4000) begin
         regblock_r_addr = rab_lite.ar_addr;
      end
      if (rab_lite.r_valid == 1 && rab_lite.ar_addr < 32'h4000) begin
         $display("Register Read detected at monitor. Address = %h, data = %h%h%h%h",regblock_r_addr,rab_lite.r_data[31:24],rab_lite.r_data[23:16],rab_lite.r_data[15:8],rab_lite.r_data[7:0]);
         if (regblock[regblock_r_addr/4] != rab_lite.r_data) begin
            $error("ERROR: Read data not correct");
            //error_num+=1;
         end
      end
   end // always_comb begin



   //////// L2 RAM Model
   //Write data to L2 model
   always_comb begin
      if (rab_lite.aw_valid == 1 && rab_lite.aw_addr >= 32'h4000) begin
         ram_addr = (rab_lite.aw_addr - 32'h4000)/4;
         if (ram_addr < 1024) begin
            va_block[ram_addr] = rab_lite.w_data;
         end else if (ram_addr < 2048) begin
            pa_block[ram_addr-1024] = rab_lite.w_data;
         end
      end
   end



   ////////////////////////////////////////////////////////////////////////////////////////
   /////////////////////////// Check axi transactions /////////////////////////////////////
   ////////////////////////////////////////////////////////////////////////////////////////
   logic [BUFFER_ADDR_BITS-1:0] addr_ptr=0, addr_check_ptr=0, aw_addr_ptr=0, aw_addr_check_ptr=0, ar_addr_ptr=0, ar_addr_check_ptr=0; // Input Buffer ptr - AW, AR channels
   logic [BUFFER_ADDR_BITS-1:0] l1_ptr=0, l1_check_ptr=0;      // L1 buffer ptr- AW, AR channels - Store if L1 hit
   logic [BUFFER_ADDR_BITS-1:0] l2_ptr=0, l2_check_ptr=0 ;     // L2 buffer ptr - AW, AR channels - Store if L1 miss
   logic [BUFFER_ADDR_BITS-1:0] out_ptr=0, out_check_ptr=0;    // Output Ordering buffer ptr - Stores order of L1, L2 transactions at output. This order will be compared with the order of data in W channel.

   // Buffers
   // axi_*_in[] -> Input Buffer
   // l1_*[] -> L1 Buffer
   // l2_*[] -> L2 Buffer
   logic [31:0]                 aw_addr_in[BUFFER_SIZE], ar_addr_in[BUFFER_SIZE], axi_addr_in;
   logic [31:0]                 l1_addr_out[BUFFER_SIZE], l2_addr_out[BUFFER_SIZE], l2_addr_in[BUFFER_SIZE];
   logic [C_AXI_ID_WIDTH-1:0]   axi_id_in, aw_id_in[BUFFER_SIZE], ar_id_in[BUFFER_SIZE], l1_id[BUFFER_SIZE], l2_id[BUFFER_SIZE];
   logic [7:0]                  aw_burst_size[BUFFER_SIZE], aw_burst_len[BUFFER_SIZE], ar_burst_size[BUFFER_SIZE], ar_burst_len[BUFFER_SIZE], axi_burst_size, axi_burst_len;
   logic [1:0]                  aw_burst_type[BUFFER_SIZE], ar_burst_type[BUFFER_SIZE], axi_burst_type;
   logic                        aw_is_write[BUFFER_SIZE], ar_is_write[BUFFER_SIZE], axi_is_write, l1_is_write[BUFFER_SIZE], l2_is_write[BUFFER_SIZE], l2_is_hit[BUFFER_SIZE], l2_is_multi[BUFFER_SIZE], l2_is_prot[BUFFER_SIZE];
   logic                        l1_multi[BUFFER_SIZE], l1_prot[BUFFER_SIZE];
   int                          out_order[BUFFER_SIZE];
   logic                        l2_is_acp[BUFFER_SIZE];
   logic                        l2_acp_saved;

   logic [31:0]                 rab_addr_in, rab_addr_in_max, exp_axi_addr_out;
   logic                        clr_rab_out; // clear L1 outputs
   logic                        exp_prot, exp_miss, exp_multi_hit, exp_acp; // L1 outputs
   logic                        exp_acp_saved;
   logic                        l2_prot, l2_miss, l2_multi_hit; // L2 outputs
   int                          exp_hit,l2_hit;
   int                          num_slices=48;
   logic [31:0]                 va_addr, va_block_entry;
   int                          set_num, set_start_addr;

   logic                        l1_was_hit,l2_was_hit; // Whether output transaction was a L1 hit or L2 hit. Used for debug.
   logic [31:0]                 l2_addr_out_debug, dropping_addr; // Used for debug.
   logic                        prot_debug,multi_debug;
   logic                        priority_is_write;
   int                          l1_prot_expected, l1_multi_expected;
   logic                        one_more_prot,one_more_multi;

   // Store incoming transactions in buffers
   always_ff @(posedge clk_i) begin
      // Write
      if (rst_ni == 0) begin
         aw_addr_ptr <= 0;
         ar_addr_ptr <= 0;
      end else if ((tgen2rab.aw_valid && tgen2rab.aw_ready) == '1) begin
         $display("AXI write coming in..addr=%h @%0d",tgen2rab.aw_addr,$time);
         aw_addr_in[aw_addr_ptr[2:0]]    <= tgen2rab.aw_addr;
         aw_id_in[aw_addr_ptr[2:0]]      <= tgen2rab.aw_id;
         aw_is_write[aw_addr_ptr[2:0]]   <= '1;
         aw_burst_size[aw_addr_ptr[2:0]] <= tgen2rab.aw_size;
         aw_burst_len[aw_addr_ptr[2:0]]  <= tgen2rab.aw_len;
         aw_burst_type[aw_addr_ptr[2:0]] <= tgen2rab.aw_burst;
         aw_addr_ptr <= aw_addr_ptr + 1'b1 ;
      end else
      //Read
      if ((tgen2rab.ar_valid && tgen2rab.ar_ready) == '1) begin
         $display("AXI read coming in..addr=%h @%0d",tgen2rab.ar_addr,$time);
         ar_addr_in[ar_addr_ptr[2:0]]    <= tgen2rab.ar_addr;
         ar_id_in[ar_addr_ptr[2:0]]      <= tgen2rab.ar_id;
         ar_is_write[ar_addr_ptr[2:0]]   <= '0;
         ar_burst_size[ar_addr_ptr[2:0]] <= tgen2rab.ar_size;
         ar_burst_len[ar_addr_ptr[2:0]]  <= tgen2rab.ar_len;
         ar_burst_type[ar_addr_ptr[2:0]] <= tgen2rab.ar_burst;
         ar_addr_ptr <= ar_addr_ptr + 1'b1;
      end
   end // always_ff @ (posedge clk_i)




/////// RAB Model /////

   // L1 TLB model
   always_comb begin
      if(aw_addr_ptr != aw_addr_check_ptr || ar_addr_ptr != ar_addr_check_ptr) begin
         // Select Read or Write based on priority if both read and write are available, else select whichever is available
         if (aw_addr_ptr != aw_addr_check_ptr && ar_addr_ptr != ar_addr_check_ptr) begin
            if (priority_is_write) begin
               axi_addr_in    = aw_addr_in[aw_addr_check_ptr[2:0]];
               axi_id_in      = aw_id_in[aw_addr_check_ptr[2:0]] ;
               axi_is_write   = aw_is_write[aw_addr_check_ptr[2:0]];
               axi_burst_size = aw_burst_size[aw_addr_check_ptr[2:0]] ;
               axi_burst_len  = aw_burst_len[aw_addr_check_ptr[2:0]] ;
               axi_burst_type = aw_burst_type[aw_addr_check_ptr[2:0]] ;
            end else begin
               axi_addr_in    = ar_addr_in[ar_addr_check_ptr[2:0]];
               axi_id_in      = ar_id_in[ar_addr_check_ptr[2:0]] ;
               axi_is_write   = ar_is_write[ar_addr_check_ptr[2:0]];
               axi_burst_size = ar_burst_size[ar_addr_check_ptr[2:0]] ;
               axi_burst_len  = ar_burst_len[ar_addr_check_ptr[2:0]] ;
               axi_burst_type = ar_burst_type[ar_addr_check_ptr[2:0]] ;
            end // else: !if(priority_is_write)
         end else if (aw_addr_ptr != aw_addr_check_ptr) begin
            axi_addr_in    = aw_addr_in[aw_addr_check_ptr[2:0]];
            axi_id_in      = aw_id_in[aw_addr_check_ptr[2:0]] ;
            axi_is_write   = aw_is_write[aw_addr_check_ptr[2:0]];
            axi_burst_size = aw_burst_size[aw_addr_check_ptr[2:0]] ;
            axi_burst_len  = aw_burst_len[aw_addr_check_ptr[2:0]] ;
            axi_burst_type = aw_burst_type[aw_addr_check_ptr[2:0]] ;
         end else if (ar_addr_ptr != ar_addr_check_ptr) begin
            axi_addr_in    = ar_addr_in[ar_addr_check_ptr[2:0]];
            axi_id_in      = ar_id_in[ar_addr_check_ptr[2:0]] ;
            axi_is_write   = ar_is_write[ar_addr_check_ptr[2:0]];
            axi_burst_size = ar_burst_size[ar_addr_check_ptr[2:0]] ;
            axi_burst_len  = ar_burst_len[ar_addr_check_ptr[2:0]] ;
            axi_burst_type = ar_burst_type[ar_addr_check_ptr[2:0]] ;
         end

         exp_axi_addr_out = 0;
         exp_hit = 0;
         rab_addr_in = axi_addr_in;
         exp_acp = 0;
         exp_acp_saved = 0;

         if(axi_burst_type==2'b01) begin // INCR burst
            rab_addr_in_max = axi_addr_in + ((axi_burst_len+1)*(1<<axi_burst_size)) - 1;
         end else begin //assume FIXED
            rab_addr_in_max = axi_addr_in + 3;
         end

         for(int i=1; i<num_slices+1; i++) begin
            if(regblock[i*8+6][0] == '1) begin // if slice is enabled
               if( (rab_addr_in >= regblock[i*8]) && (rab_addr_in_max < regblock[i*8+2]) ) begin // hit
                  if (exp_hit == 0) begin // In case of 2 hits, out addr is addr in first slice
                     exp_axi_addr_out = regblock[i*8+4] + rab_addr_in - regblock[i*8];
                  end
                  exp_hit+=1;
                  if ((regblock[i*8+6][2] == '0 && axi_is_write == '1) || (regblock[i*8+6][1] == '0 && axi_is_write == '0)) begin // if protected
                     exp_prot = 1;
                     exp_axi_addr_out = rab_addr_in;
                  end else begin
                     exp_prot = 0;
                  end
                  if (regblock[i*8+6][3] == '1) begin
                     exp_acp_saved = '1;
                  end
               end
            end // if (regblock[i*4+3][0] == '1)
         end // for (int i=1; i<num_slices+1; 1++)

         if(exp_hit > 2) begin // multi_hit
            exp_multi_hit = '1;
            exp_miss = '0;
         end else if (exp_hit == 0) begin // miss
            exp_miss = '1;
            exp_multi_hit = '0;
         end else begin // hit
            exp_miss = '0;
            exp_multi_hit = '0;
         end
         if (exp_prot ==0 && exp_multi_hit ==0 && exp_miss==0) begin
            exp_acp = exp_acp_saved;
         end
      end // if (addr_ptr != addr_check_ptr)
      else if (clr_rab_out) begin
         exp_prot = '0;
         exp_hit = 0;
         exp_miss = '0;
         exp_multi_hit = '0;
         exp_acp = '0;
         exp_acp_saved = '0;
      end
   end // always_comb begin

   // Move transaction to L1/L2 buffer based on L1 TLB output.
   // L1 buffer => L1 Hit
   // L2 buffer => L1 Miss

   always_ff @(posedge clk_i) begin
      if (rst_ni == 0) begin
         priority_is_write <= 0;
      end else if(exp_miss) begin
         l2_addr_in[l2_ptr[2:0]]  <= axi_addr_in;
         l2_is_write[l2_ptr[2:0]] <= axi_is_write;
         l2_id[l2_ptr[2:0]]       <= axi_id_in;
         l2_ptr                   <= l2_ptr + 1'b1;
         clr_rab_out <= 1;
         if (axi_is_write) begin
            aw_addr_check_ptr           <= aw_addr_check_ptr + 1'b1;
            priority_is_write <= 1;
         end else begin
            ar_addr_check_ptr           <= ar_addr_check_ptr + 1'b1;
            priority_is_write <= 0;
         end
      end else if (exp_hit>0 && exp_acp==0) begin
         l1_addr_out[l1_ptr[2:0]] <= exp_axi_addr_out;
         l1_is_write[l1_ptr[2:0]] <= axi_is_write;
         l1_id[l1_ptr[2:0]]       <= axi_id_in;
         l1_prot[l1_ptr[2:0]]     <= exp_prot;
         l1_multi[l1_ptr[2:0]]    <= exp_multi_hit;
         l1_ptr                   <= l1_ptr + 1'b1;
         clr_rab_out <= 1;
         if (axi_is_write) begin
            aw_addr_check_ptr           <= aw_addr_check_ptr + 1'b1;
            priority_is_write <= 1;
         end else begin
            ar_addr_check_ptr           <= ar_addr_check_ptr + 1'b1;
            priority_is_write <= 0;
         end
      end else if (exp_acp) begin // if (exp_hit>0 && exp_axp==0)
         clr_rab_out <= 1;
         if (axi_is_write) begin
            aw_addr_check_ptr           <= aw_addr_check_ptr + 1'b1;
            priority_is_write <= 1;
         end else begin
            ar_addr_check_ptr           <= ar_addr_check_ptr + 1'b1;
            priority_is_write <= 0;
         end
      end else begin
         clr_rab_out <= 1;
      end // else: !if(exp_hit>0)
      l1_prot_expected <= exp_prot;
      l1_multi_expected <= exp_multi_hit;
   end // always_ff @ (clk_i)

   ///// L2 TLB model
   // Check L2 TLB for hit/miss
   always_comb begin
      if (l2_ptr != l2_check_ptr) begin
         l2_hit = 0;
         l2_prot = 0;
         l2_multi_hit = 0;
         l2_miss = 0;
         l2_acp_saved = 0;
         va_addr = l2_addr_in[l2_check_ptr[2:0]];
         set_num = va_addr[12+5-1:12]; // 32 sets, Page size = 4k. TODO: Parameterise
         set_start_addr = set_num * 16*2; // TODO: Parameterise
         for(int j=0; j<32; j++) begin //16*2 entries in set. TODO: Parameterise
            va_block_entry = va_block[set_start_addr+j];
            if((va_addr[31:12] == va_block_entry[23:4]) && va_block_entry[0]) begin // L2 hit
               l2_hit+=1;
               if ((l2_is_write[l2_check_ptr[2:0]] && ~va_block_entry[2]) || (~l2_is_write[l2_check_ptr[2:0]] && ~va_block_entry[1])) begin //prot
                  l2_prot = 1;
               end else begin
                  if(l2_hit == 1) begin
                     l2_addr_out[l2_check_ptr[2:0]] = {pa_block[set_start_addr+j][19:0],l2_addr_in[l2_check_ptr[2:0]][11:0]};
                     l2_addr_out_debug = {pa_block[set_start_addr+j][19:0],l2_addr_in[l2_check_ptr[2:0]][11:0]};
                  end
               end
               l2_acp_saved = va_block_entry[3];
            end
         end // for (int j=0; j<16; j++)
         if(l2_hit == 0) begin
            l2_miss = 1;
         end else if (l2_hit > 1) begin
            l2_miss = 0;
`ifdef TLB_MULTIHIT
            l2_multi_hit = 1;
`endif
         end else begin
            l2_miss = 0;
         end

         l2_is_hit[l2_check_ptr[2:0]] = ~l2_miss;
         l2_is_multi[l2_check_ptr[2:0]] = l2_multi_hit;
         l2_is_prot[l2_check_ptr[2:0]] = l2_prot;
         l2_is_acp[l2_check_ptr[2:0]] = l2_acp_saved && ~l2_multi_hit;
      end
   end // always_comb begin
///////////////////

   /// RAB Output transactions
   logic [C_AXI_ID_WIDTH-1:0]   aw_id_out,ar_id_out;
   logic                        axi_out_is_write;
   logic [31:0]                 aw_addr_out, ar_addr_out ;

   always_comb begin
      if((rab2mem.aw_valid && rab2mem.aw_ready) == 1) begin // Write
         aw_addr_out = rab2mem.aw_addr;
         aw_id_out = rab2mem.aw_id;
//         axi_out_is_write = 1;
      end
      if((rab2mem.ar_valid && rab2mem.ar_ready) == 1) begin //Read
         ar_addr_out <= rab2mem.ar_addr;
         ar_id_out <= rab2mem.ar_id;
//         axi_out_is_write = 0;
      end
   end

   logic    intr_miss_o_d, intr_prot_o_d, intr_multi_o_d;
   int      p_debug = 0;
   /// Compare AXI AW, AR outputs with those in Buffers
   always_ff @(posedge clk_i) begin
      //Write
      if ((rab2mem.aw_valid && rab2mem.aw_ready) == 1) begin
         if ((aw_id_out == l1_id[l1_check_ptr[2:0]]) && (aw_addr_out == l1_addr_out[l1_check_ptr[2:0]]) && (l1_is_write[l1_check_ptr[2:0]]==1) && l1_check_ptr != l1_ptr)begin
            $display("L1 Hit!! AXI write going out..addr = %h",aw_addr_out);
            l1_check_ptr <= l1_check_ptr + 1'b1;
//            l1_was_hit <= 1;
//            l2_was_hit <= 0;
            out_order[out_ptr[2:0]] <= 1;
            out_ptr <= out_ptr + 1'b1;
         end else if ((aw_id_out == l2_id[l2_check_ptr[2:0]]) && (aw_addr_out == l2_addr_out[l2_check_ptr[2:0]]) && (l2_is_write[l2_check_ptr[2:0]]==1) && l2_check_ptr != l2_ptr) begin
            $display("L2 Hit!! AXI write going out..addr = %h",aw_addr_out);
            if (l2_is_hit[l2_check_ptr[2:0]] == 0) begin
               $error("Expected Miss");
               error_miss+=1;
            end
            l2_check_ptr <= l2_check_ptr + 1'b1;
            l1_was_hit <= 0;
            l2_was_hit <= 1;
            out_order[out_ptr[2:0]] <= 2;
            out_ptr <= out_ptr + 1'b1;
         end else begin
            $error("Unexpected AXI write going out. AXI Addr = %h, AXI ID = %h, time=%t",aw_addr_out,aw_id_out,$time);
            //$display("aw_id_out = %h, l1_id = %h, l2_id = %h", aw_id_out, l1_id[l1_check_ptr[2:0]], l2_id[l2_check_ptr[2:0]]);
            error_axi+=1;
//            l1_was_hit <= 0;
//            l2_was_hit <= 0;
         end // else: !if((aw_id_out == l2_id[l2_check_ptr[2:0]]) && (aw_addr_out == l2_addr_out[l2_check_ptr[2:0]]) && (l2_is_write[l2_check_ptr[2:0]]==1) && l2_check_ptr != l2_ptr)
         // if a miss, prot or multi is seen at the output along with a valid write transaction.
         intr_miss_o_d <= intr_miss_o && (l2_ptr != l2_check_ptr && ~l2_is_hit[l2_check_ptr[2:0]]) && l2_is_write[l2_check_ptr[2:0]];
         intr_prot_o_d <= intr_prot_o && (l2_ptr != l2_check_ptr && l2_is_prot[l2_check_ptr[2:0]]) && l2_is_write[l2_check_ptr[2:0]];
         intr_multi_o_d <= intr_multi_o && (l2_ptr != l2_check_ptr && l2_is_multi[l2_check_ptr[2:0]]) && l2_is_write[l2_check_ptr[2:0]];
      end else if (((intr_miss_o && (l2_check_ptr != l2_ptr) && l2_is_write[l2_check_ptr[2:0]])|| intr_miss_o_d)) begin
         out_order[out_ptr[2:0]] <= 0;
         out_ptr <= out_ptr + 1'b1;
         dropping_addr <= l2_addr_in[l2_check_ptr[2:0]];
         intr_miss_o_d <= 0;
      end else if ( ((intr_prot_o && (l2_check_ptr != l2_ptr)) && ~one_more_prot && l2_is_prot[l2_check_ptr[2:0]] && l2_is_write[l2_check_ptr[2:0]])||intr_prot_o_d) begin
         out_order[out_ptr[2:0]] <= 10;
         out_ptr <= out_ptr + 1'b1;
         dropping_addr <= l2_addr_in[l2_check_ptr[2:0]];
         intr_prot_o_d <= 0;
         p_debug <= p_debug + 1;
      end else if ( ((intr_multi_o && (l2_check_ptr != l2_ptr)) && ~one_more_multi && l2_is_multi[l2_check_ptr[2:0]] && l2_is_write[l2_check_ptr[2:0]])||intr_multi_o_d) begin
         out_order[out_ptr[2:0]] <= 20;
         out_ptr <= out_ptr + 1'b1;
         dropping_addr <= l2_addr_in[l2_check_ptr[2:0]];
         intr_multi_o_d <= 0;
      end else if(l2_is_acp[l2_check_ptr[2:0]] && (l2_check_ptr != l2_ptr) && l2_is_write[l2_check_ptr[2:0]]) begin
         l2_check_ptr <= l2_check_ptr + 1'b1;
         out_order[out_ptr[2:0]] <= 30;
         out_ptr <= out_ptr + 1'b1;
      end else if(l2_is_acp[l2_check_ptr[2:0]] && (l2_check_ptr != l2_ptr) && ~l2_is_write[l2_check_ptr[2:0]]) begin
         l2_check_ptr <= l2_check_ptr + 1'b1;
      end
      // out_order is used to keep track of write transaction results. It will be used to validate/drop the W channel signals.

      //Read
      if ((rab2mem.ar_valid && rab2mem.ar_ready) == 1) begin
         if ((ar_id_out == l1_id[l1_check_ptr[2:0]]) && (ar_addr_out == l1_addr_out[l1_check_ptr[2:0]]) && (l1_is_write[l1_check_ptr[2:0]]==0) && l1_check_ptr != l1_ptr) begin
            $display("L1 Hit!! AXI read going out..addr = %h",ar_addr_out);
            l1_check_ptr <= l1_check_ptr + 1'b1;
         end else if ((ar_id_out == l2_id[l2_check_ptr[2:0]]) && (ar_addr_out == l2_addr_out[l2_check_ptr[2:0]]) && (l2_is_write[l2_check_ptr[2:0]]==0) && l2_check_ptr != l2_ptr) begin
            $display("L2 Hit!! AXI read going out..addr = %h",ar_addr_out);
            l2_check_ptr <= l2_check_ptr + 1'b1;
         end else begin
            $error("Unexpected AXI read going out. AXI Addr = %h, AXI ID = %h, time=%t",ar_addr_out,ar_id_out,$time);
            error_axi+=1;
         end
      end // if ((rab2mem.ar_valid && rab2mem.ar_ready) == 1)


   end



   ////////////// Write Channel //////////////////////////////////
   logic [6:0]                 w_ptr=0, w_check_ptr=0; // Ptr - Input buffer
   logic [6:0]                 hit_ptr=0,hit_check_ptr=0; // Ptr - Used to store order of L1 Hit and Miss.
   logic [6:0]                 l1_w_ptr=0,l2_w_ptr=0,l1_w_check_ptr=0,l2_w_check_ptr=0; // Ptr - L1 and L2 buffer
   //Buffers
   logic [63:0]                wdata[64],l1_wdata[64],l2_wdata[64],l2_wdata_debug,l1_wdata_debug,dropping_data;
   logic                       wlast[64],l1_wlast[64],l2_wlast[64];
   int                         l1_hit[64]; // Store if L1 hit or L1 miss or L1 multi/prot.

   logic                       waiting_last_drop, second_miss;
   logic                       wlast_received;
   int                         error_wdata=0;
   logic                       debug_signal,input_debug; // Used for Debug
   int                         out_debug; // Used for Debug
   logic [31:0]                wdebug_addr[64], current_addr_debug; // Used for Debug

   logic [BUFFER_ADDR_BITS-1:0]                 l2_wlast_ptr=0, l2_wlast_check_ptr=0;
   logic [6:0]                                  wlast_idx[BUFFER_SIZE];

   // Store inputs in In buffer
   always_ff @(posedge clk_i) begin
      if (rst_ni == 0) begin
         w_ptr <= 0;
      end else if ((tgen2rab.w_valid && tgen2rab.w_ready) == '1) begin
         wdata[w_ptr[5:0]] <= tgen2rab.w_data;
         wlast[w_ptr[5:0]] <= tgen2rab.w_last;
         w_ptr <= w_ptr + 1'b1;
      end
   end

   // Store RAB hit/miss. To be used for W channel
   always_ff @(posedge clk_i) begin
      if((exp_miss) && axi_is_write) begin
         l1_hit[hit_ptr[5:0]] <= 0;
         wdebug_addr[hit_ptr[5:0]] <= axi_addr_in;
         hit_ptr <= hit_ptr + 1'b1;
      end else if ( (exp_prot || exp_multi_hit || exp_acp) && axi_is_write) begin
         l1_hit[hit_ptr[5:0]] <= 2;
         hit_ptr <= hit_ptr + 1'b1;
      end else if (exp_hit>0 && axi_is_write) begin
         l1_hit[hit_ptr[5:0]] <= 1;
         wdebug_addr[hit_ptr[5:0]] <= exp_axi_addr_out;
         hit_ptr <= hit_ptr + 1'b1;
      end
   end // always_ff @ (posedge clk_i)

   logic [6:0] debug_wlast_idx;
   // Move w channel signals from In buffer to L1/L2 buffers. Do not move if In buffer is empty.
   always_ff @(posedge clk_i) begin
      if(l1_hit[hit_check_ptr[5:0]] == 0 && hit_check_ptr != hit_ptr && w_check_ptr != w_ptr) begin // L1 miss/prot/multi. Move to L2 Buffer.
         l2_wdata[l2_w_ptr[5:0]]  <= wdata[w_check_ptr[5:0]];
         l2_wlast[l2_w_ptr[5:0]]  <= wlast[w_check_ptr[5:0]];
         w_check_ptr              <= w_check_ptr + 1'b1;
         l2_w_ptr                 <= l2_w_ptr + 1'b1;
         l2_wdata_debug  <= wdata[w_check_ptr[5:0]];
         input_debug <= wlast[w_check_ptr[5:0]];
         current_addr_debug <= wdebug_addr[hit_check_ptr[5:0]];
         if(wlast[w_check_ptr[5:0]]) begin
            hit_check_ptr <= hit_check_ptr + 1'b1;
            wlast_idx[l2_wlast_ptr[2:0]] <= l2_w_ptr;
            debug_wlast_idx <= l2_w_ptr;
            l2_wlast_ptr <= l2_wlast_ptr + 1'b1;
         end
      end else if (l1_hit[hit_check_ptr[5:0]] == 1 && hit_check_ptr != hit_ptr && w_check_ptr != w_ptr) begin // L1 hit. Move to L1 Buffer.
         l1_wdata[l1_w_ptr[5:0]]  <= wdata[w_check_ptr[5:0]];
         l1_wlast[l1_w_ptr[5:0]]  <= wlast[w_check_ptr[5:0]];
         w_check_ptr              <= w_check_ptr + 1'b1;
         l1_w_ptr                 <= l1_w_ptr + 1'b1;
         l1_wdata_debug  <= wdata[w_check_ptr[5:0]];
         current_addr_debug <= wdebug_addr[hit_check_ptr[5:0]];
         if(wlast[w_check_ptr[5:0]])
           hit_check_ptr <= hit_check_ptr + 1'b1;
      end else if (l1_hit[hit_check_ptr[5:0]] == 2 && hit_check_ptr != hit_ptr && w_check_ptr != w_ptr) begin // L1 multi/prot. Drop data.
         w_check_ptr              <= w_check_ptr + 1'b1;
         if(wlast[w_check_ptr[5:0]])
           hit_check_ptr <= hit_check_ptr + 1'b1;
      end
   end // always_ff @ (clk_i)



   logic check_now, waiting_wlast;
   assign check_now = rab2mem.w_valid && rab2mem.w_ready && rab2mem.aw_valid && rab2mem.aw_ready;
   always_ff @(posedge clk_i) begin
      if (rst_ni == 0) begin
         waiting_wlast <= 0;
      end else if (rab2mem.w_valid && rab2mem.w_ready) begin
         waiting_wlast <= ~rab2mem.w_last;
      end
   end

   // compare w channel signals
   always_ff @(posedge clk_i) begin
      if(((out_order[out_check_ptr[2:0]]==1 && out_check_ptr != out_ptr)||(check_now&&~waiting_wlast&&out_check_ptr == out_ptr)) && (wlast_received || l1_w_check_ptr != l1_w_ptr)) begin // This was a L1 hit
         if(wlast_received) begin
            wlast_received <= 0;
            out_check_ptr <= out_check_ptr + 1'b1;
         end
         if((rab2mem.w_valid && rab2mem.w_ready) == '1) begin  // valid wdata
            if(rab2mem.w_data == l1_wdata[l1_w_check_ptr[5:0]]) begin
               $display("L1.wdata correct. wdata = %h, time=%t",l1_wdata[l1_w_check_ptr[5:0]],$time);
               l1_w_check_ptr <= l1_w_check_ptr + 1'b1;
               if(rab2mem.w_last == 1 && l1_wlast[l1_w_check_ptr[5:0]] == 1) begin // wlast. Trans completed.
                  out_check_ptr <= out_check_ptr + 1'b1;
               end
            end else begin
               $error("wdata not correct.L1. Expected = %h, Actual = %h, time=%t",l1_wdata[l1_w_check_ptr[5:0]],rab2mem.w_data,$time);
               error_wdata+=1;
               l1_w_check_ptr <= l1_w_check_ptr + 1'b1;
            end
         end
      end else if(out_order[out_check_ptr[2:0]]==2 && out_check_ptr != out_ptr && l2_w_ptr != l2_w_check_ptr) begin // This was L2 hit
         if((rab2mem.w_valid && rab2mem.w_ready) == '1) begin // valid wdata
            if(rab2mem.w_data == l2_wdata[l2_w_check_ptr[5:0]]) begin
               $display("L2.wdata correct. wdata = %h",l2_wdata[l2_w_check_ptr[5:0]]);
               l2_w_check_ptr <= l2_w_check_ptr + 1'b1;
               if(rab2mem.w_last == 1 && l2_wlast[l2_w_check_ptr[5:0]] == 1) begin // wlast. Trans completed.
                  out_check_ptr <= out_check_ptr + 1'b1;
                  l2_wlast_check_ptr <= l2_wlast_check_ptr + 1'b1;
               end
            end else begin
               $error("wdata not correct.L2. Expected = %h, Actual = %h, time=%t",l2_wdata[l2_w_check_ptr[5:0]],rab2mem.w_data,$time);
               error_wdata+=1;
               l2_w_check_ptr <= l2_w_check_ptr + 1'b1;
            end
         end
      end else if (out_order[out_check_ptr[2:0]]%10==0 && out_check_ptr != out_ptr && l2_w_ptr != l2_w_check_ptr) begin // L2 miss. Drop w channel signals.
         //if(intr_miss_o || intr_multi_o || intr_prot_o || waiting_last_drop) begin
         if (l2_wlast_check_ptr != l2_wlast_ptr) begin
            l2_w_check_ptr <= wlast_idx[l2_wlast_check_ptr[2:0]];
         end else begin
            l2_w_check_ptr <= l2_w_check_ptr + 1'b1;
         end
         dropping_data <= l2_wdata[l2_w_check_ptr[5:0]];
         if (l2_wlast[l2_w_check_ptr[5:0]]) begin
            out_check_ptr <= out_check_ptr + 1'b1;
            l2_wlast_check_ptr <= l2_wlast_check_ptr + 1'b1;
            l2_w_check_ptr <= l2_w_check_ptr + 1'b1;
         end
         if( (rab2mem.w_valid && rab2mem.w_ready) == '1) begin // wdata received for L1 Hit when dropping data
            if(rab2mem.w_data == l1_wdata[l1_w_check_ptr[5:0]]) begin
               $display("L1.wdata correct. wdata = %h",l1_wdata[l1_w_check_ptr[5:0]]);
               l1_w_check_ptr <= l1_w_check_ptr + 1'b1;
            end else begin
               $error("wdata not correct.L1. Expected = %h, Actual = %h, time=%t",l1_wdata[l1_w_check_ptr[5:0]],rab2mem.w_data,$time);
               error_wdata+=1;
               l1_w_check_ptr <= l1_w_check_ptr + 1'b1;
            end
            if (rab2mem.w_last == 1) begin
               wlast_received <= 1;
            end
         end
         //end
      end

      debug_signal <= l2_wlast[l2_w_check_ptr[5:0]];
      out_debug <= out_order[out_check_ptr[2:0]];

   end // always_ff @ (posedge clk_i)


   //////////////////////////////////////////////////////////////////////////////////
   /////////////////// Check miss, multi, prot //////////////////////////////////////
   //////////////////////////////////////////////////////////////////////////////////
   logic [31:0] l1_check_addr, l2_check_addr;
   always_ff @(posedge clk_i) begin
      if (rst_ni == 0) begin
         one_more_prot <= 0;
         one_more_multi <= 0;
      end else
      if(intr_miss_o) begin
         if(l2_ptr != l2_check_ptr && l2_is_hit[l2_check_ptr[2:0]]) begin
            $error("Unexpected Miss, time=%t",$time);
            error_miss+=1;
            l2_check_ptr <= l2_check_ptr + 1'b1;
         end else if (l2_ptr != l2_check_ptr && ~l2_is_hit[l2_check_ptr[2:0]])begin
            $display("L2 Miss!! addr = %h, ID = %h, time=%t",l2_addr_in[l2_check_ptr[2:0]],l2_id[l2_check_ptr[2:0]],$time);
            l2_check_ptr <= l2_check_ptr + 1'b1;
         end
      end //else
      if(intr_prot_o) begin
         l1_check_addr <= l1_addr_out[l1_check_ptr[2:0]];
         l2_check_addr <= l2_addr_in[l2_check_ptr[2:0]];
         if (one_more_prot == 1) begin
            one_more_prot <= 0;
            $display("Prot!! Not sure L1 or L2. Another Prot would have been detected a little earlier.");
         end else if ((l2_ptr != l2_check_ptr && l2_is_prot[l2_check_ptr[2:0]]) && (l1_ptr != l1_check_ptr && l1_prot[l1_check_ptr[2:0]])) begin
            $display("Prot!! Not sure L1 or L2. Another Prot expected soon.");
            l2_check_ptr <= l2_check_ptr + 1'b1;
            l1_check_ptr <= l1_check_ptr + 1'b1;
            one_more_prot <= 1;
         end else if (l2_ptr != l2_check_ptr && l2_is_prot[l2_check_ptr[2:0]]) begin
            $display("L2.Prot!! addr = %h, ID = %h, RW_type=%d",l2_addr_in[l2_check_ptr[2:0]],l2_id[l2_check_ptr[2:0]],l2_is_write[l2_check_ptr[2:0]]);
            l2_check_ptr <= l2_check_ptr + 1'b1;
         end else if (l1_ptr != l1_check_ptr && l1_prot[l1_check_ptr[2:0]]) begin
            $display("L1.Prot!!addr = %h, ID = %h, RW_type=%d, time=%t",l1_addr_out[l1_check_ptr[2:0]],l1_id[l1_check_ptr[2:0]],l1_is_write[l1_check_ptr[2:0]],$time);
            l1_check_ptr <= l1_check_ptr + 1'b1;
         end else begin
            $error("Unexpected Prot, time=%t",$time);
            error_miss+=1;
         end
      end //else
      if(intr_multi_o) begin
         if (one_more_multi == 1) begin
            one_more_multi <= 0;
            $display("Multi!! Not sure L1 or L2. Another Multi would have been detected a little earlier.");
         end else if ((l2_ptr != l2_check_ptr && l2_is_multi[l2_check_ptr[2:0]]) && (l1_ptr != l1_check_ptr && l1_multi[l1_check_ptr[2:0]])) begin
            $display("Multi!! Not sure L1 or L2. Another Multi expected soon.");
            l2_check_ptr <= l2_check_ptr + 1'b1;
            l1_check_ptr <= l1_check_ptr + 1'b1;
            one_more_multi <= 1;
         end else if (l2_ptr != l2_check_ptr && l2_is_multi[l2_check_ptr[2:0]]) begin
            $display("L2.Multi!! addr = %h, ID = %h, RW_type=%d",l2_addr_in[l2_check_ptr[2:0]],l2_id[l2_check_ptr[2:0]],l2_is_write[l2_check_ptr[2:0]]);
            l2_check_ptr <= l2_check_ptr + 1'b1;
         end else if (l1_ptr != l1_check_ptr && l1_multi[l1_check_ptr[2:0]]) begin
            $display("L1.Multi!!ID = %h, RW_type=%d",l1_id[l1_check_ptr[2:0]],l1_is_write[l1_check_ptr[2:0]]);
            l1_check_ptr <= l1_check_ptr + 1'b1;
         end else begin
            $error("Unexpected Multi, time=%t",$time);
            error_miss+=1;
         end
      end
   end // always_ff @ (posedge clk_i)
   // one_more_multi and one_more_prot are required because we cannot distinguish between the multi/prot generated from L1 TLB and L2 TLB at RAB output.
   // If we expect a multi/prot from both L1 and L2, we assert these signals and make sure another multi/prot is detected.


   /// Number of errors
   always_comb begin
      error_num = error_axi + error_miss + error_buf + error_wdata;
   end
//




endmodule
